// NOTES:
// Not sure what to output

module score ( input         Clk,                // 50 MHz clock
                             Reset_Score,        // Active-high reset signal
                             frame_clk,          // The clock indicating a new frame (~60Hz)
									  
					input logic collision_blue, collision_red,
               output logic 
);

endmodule